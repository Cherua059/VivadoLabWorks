`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.02.2025 15:02:07
// Design Name: 
// Module Name: shifter_32_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module shifter_32_tb();

    reg [31 : 0] a;
    reg [4 : 0] b;
    reg [1 : 0] c;
    wire [31 : 0] z;
    
    shifter_32 shift32 (.a(a), .b(b), .c(c), .z(z));
    
    initial
        begin
        $monitor("Input = %b, Shift Amount = %b, Shift type = %b, Output = %b", a, b, c, z);
        
            a = 32'b01111111111111111111111111111111; b = 5'b00000; c = 2'b01; //no shift
        
        #50 a = 32'b11111111111111111111111111111111; b = 5'b10000; c = 2'b01; //(or) c = 2'b00 //16 BIT LS
        #50 a = 32'b11111111111111111111111111111111; b = 5'b10000; c = 2'b11; //16 BIT ARS
        #50 a = 32'b11111111111111111111111111111111; b = 5'b10000; c = 2'b10; //16 BIT LRS
        
        #50 a = 32'b01111111111111111111111111111111; b = 5'b01000; c = 2'b01; //(or) c = 2'b00 //8 BIT LS
        #50 a = 32'b01111111111111111111111111111111; b = 5'b01000; c = 2'b11; //8 BIT ARS
        #50 a = 32'b01111111111111111111111111111111; b = 5'b01000; c = 2'b10; //8 BIT LRS
        
        #50 a = 32'b11111111111111111111111111111111; b = 5'b00100; c = 2'b01; //(or) c = 2'b00 //4 BIT LS
        #50 a = 32'b11111111111111111111111111111111; b = 5'b00100; c = 2'b11; //4 BIT ARS
        #50 a = 32'b11111111111111111111111111111111; b = 5'b00100; c = 2'b10; //4 BIT LRS
        
        #50 a = 32'b01111111111111111111111111111111; b = 5'b00010; c = 2'b01; //(or) c = 2'b00 //2 BIT LS
        #50 a = 32'b01111111111111111111111111111111; b = 5'b00010; c = 2'b11; //2 BIT ARS
        #50 a = 32'b01111111111111111111111111111111; b = 5'b00010; c = 2'b10; //2 BIT LRS
        
        #50 a = 32'b11111111111111111111111111111111; b = 5'b00001; c = 2'b01; //(or) c = 2'b00 //1 BIT LS
        #50 a = 32'b11111111111111111111111111111111; b = 5'b00001; c = 2'b11; //1 BIT ARS
        #50 a = 32'b11111111111111111111111111111111; b = 5'b00001; c = 2'b10; //1 BIT LRS
        
        #50 a = 32'b01111111111111111111111111111111; b = 5'b11111; c = 2'b01; //(or) c = 2'b00 //32 BIT LS
        #50 a = 32'b01111111111111111111111111111111; b = 5'b11111; c = 2'b11; //32 BIT ARS
        #50 a = 32'b01111111111111111111111111111111; b = 5'b11111; c = 2'b10; //32 BIT LRS
        $finish;
        end

endmodule
